`ifndef CYCLE
	`define CYCLE 10
`endif

`ifndef Tdrive
	`define Tdrive #(2)
`endif

`timescale 1ns/1ns
