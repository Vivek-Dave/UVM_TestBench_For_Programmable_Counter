
`include "interface.sv"
`include "tb_pkg.sv"
module top;
  import uvm_pkg::*;
  import tb_pkg::*;
  
  bit clk; // external signal declaration

  //----------------------------------------------------------------------------
  dut_if i_intf(clk);
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  pcnt DUT(.din(i_intf.din),
		   .dout(i_intf.dout),
		   .ld(i_intf.ld),
		   .inc(i_intf.inc),
		   .clk(i_intf.clk),
		   .rst_n(i_intf.rst_n)
          );
  //----------------------------------------------------------------------------               
  
  initial begin
    clk<=0;
  end
  
  always #5 clk=~clk;
  
  //----------------------------------------------------------------------------
  initial begin
    $dumpfile("dumpfile.vcd");
    $dumpvars;
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    uvm_config_db#(virtual dut_if)::set(uvm_root::get(),"","vif",i_intf);
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    run_test("test");
  end
  //----------------------------------------------------------------------------
endmodule

